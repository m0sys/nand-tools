module thruwire (
    // OUTPUTS
    output o_led

    // INPUTS
    ,input i_sw
    );

    assign o_led = i_sw;
endmodule
