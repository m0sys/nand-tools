// Gate-lvl desc of 4bit add-sub circuit (Fig. 4.13).

module circ_437
endmodule
