// Top module for rtl design exercise 8.7.

module rtl_design607 #(parameter WIDTH=8)  (
    // OUTPUTS
    output [WIDTH-1:0] RA_o
    ,output carry_o

    // INPUTS
    ,input start_i
    ,input clk_i
    ,input rst_b_i
    );
endmodule
